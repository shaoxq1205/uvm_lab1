/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s8a/s8adaaad896791bac-1.4-1349388157-0