/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sd8/sd820911d6a6c6a89-1.4-1349388122-0