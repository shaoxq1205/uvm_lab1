/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sbd/sbd027f2d165a2710-1.4-1349388226-0