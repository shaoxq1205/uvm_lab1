/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s8b/s8bfe92d89057018d-1.4-1349388236-0