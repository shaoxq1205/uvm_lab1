/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sfa/sfa011b16c4167145-1.4-1349388231-0