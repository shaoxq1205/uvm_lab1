/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s0d/s0de8a2eee147b57e-1.4-1349388072-0