/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s8c/s8cf9ed5cc949ce3f-1.3-1349388147-0