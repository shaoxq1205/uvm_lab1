/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s86/s865590d08c8fcb33-1.4-1349388016-0