/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sf8/sf8e12157157e6f98-1.4-1349388154-0