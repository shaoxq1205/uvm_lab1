/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sc2/sc2cf1cce1cac5411-1.4-1349388093-0