/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s00/s00873edc873f5184-1.4-1349388157-0