/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/se4/se4c52b10c2c083bd-1.4-1349388184-0