/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s6f/s6f40a6d37caa621c-1.4-1349388136-0