/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sa4/sa4c90356ebf1896d-1.3-1349388180-0