/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s91/s91f7c8e97b129490-1.4-1349387987-0