/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s9b/s9b631a733bc3f574-1.4-1349388198-0