/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sd4/sd4e6d4e67a9cf209-1.4-1349388178-0