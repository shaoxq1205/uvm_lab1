/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sf5/sf5afbcc0f42e6724-1.3-1349388148-0