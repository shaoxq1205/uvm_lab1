/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sbc/sbcf337c9235160f7-1.4-1349388089-0