/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s66/s66c4b7291b4ff2cc-1.4-1349388133-0