/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s27/s2798bf6b43873beb-1.4-1349388012-0