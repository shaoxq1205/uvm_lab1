/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sbd/sbd03c95c2e4157ee-1.4-1349388132-0