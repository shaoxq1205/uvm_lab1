/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s2b/s2b91a21664dfa6d1-1.4-1349388006-0