/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s76/s767221b61a67e75f-1.4-1349388039-0