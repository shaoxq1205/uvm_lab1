/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s81/s812eede47c570b4d-1.4-1349388162-0