/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/seb/seb025d8bbc926f15-1.4-1349388141-0