/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s65/s654172f181a4d6d7-1.4-1349387966-0