/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sd4/sd4a0c5786246564a-1.4-1349388190-0