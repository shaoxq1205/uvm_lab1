/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s73/s732a4381047161c3-1.4-1349388121-0