/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s8d/s8dca0fb15a0153a6-1.1-1300484144-0