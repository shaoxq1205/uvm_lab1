/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s0a/s0aede92fa7ee3247-1.4-1349388019-0