/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sbd/sbd2fbfdc931ac127-1.4-1349388092-0