/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sb2/sb27680b2d477075f-1.4-1349388011-0