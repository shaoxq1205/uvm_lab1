/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s9e/s9e8fb2195d5682fc-1.4-1349387993-0