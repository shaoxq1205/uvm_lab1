/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s15/s153a12bc899d1b8d-1.4-1349388197-0