/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s1b/s1bd5e4b42c15c54b-1.4-1349388152-0