/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sda/sda33e36c497c3ea8-1.5-1350508138-0