/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sb6/sb648bde2447785eb-1.4-1349388154-0