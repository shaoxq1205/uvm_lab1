/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s8a/s8ac8b6557d21d6f0-1.3-1349388146-0