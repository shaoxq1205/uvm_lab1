library verilog;
use verilog.vl_types.all;
entity pcounter_test_pkg is
end pcounter_test_pkg;
