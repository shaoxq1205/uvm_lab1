/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s81/s81f4072b72329b3f-1.4-1349388001-0