/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s52/s52ca7cb8c48c662d-1.3-1349388100-0