/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s1a/s1aca4b12e9134fc5-1.4-1349388006-0