/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sf1/sf145357a21833e7f-1.4-1349388025-0