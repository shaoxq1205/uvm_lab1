library verilog;
use verilog.vl_types.all;
entity quvm_addons_pkg is
end quvm_addons_pkg;
