/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s58/s5808692f501a23ed-1.3-1349388149-0