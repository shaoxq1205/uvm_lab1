library verilog;
use verilog.vl_types.all;
entity XlSvResetGeneratorPkg is
end XlSvResetGeneratorPkg;
