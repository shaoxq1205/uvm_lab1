/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s9f/s9f3c2dd2eb2dd89d-1.4-1349388002-0