/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s14/s144bb68490c4ec4c-1.4-1349387965-0