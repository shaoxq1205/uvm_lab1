/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s47/s47ea3133dcf99681-1.4-1349388177-0