/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s8c/s8c0b47a23dbb4b1a-1.4-1349388154-0