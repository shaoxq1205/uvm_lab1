/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s48/s480798a0ecdf699b-1.3-1349388148-0