/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sd0/sd05215b5b8930f7d-1.4-1349388021-0