/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sf0/sf07c045d904e58c8-1.4-1349387998-0