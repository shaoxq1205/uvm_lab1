/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s8a/s8a61e3898c119086-1.4-1349388038-0