/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sf4/sf46351626c6e25a3-1.4-1349387987-0