/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sc5/sc514e355dba5fafc-1.4-1349388181-0