/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s4a/s4aed3e1faf64c7eb-1.4-1349388120-0