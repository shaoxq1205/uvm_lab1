/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s27/s275daa36d5dd965a-1.4-1349388078-0