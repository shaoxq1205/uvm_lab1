/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s01/s01f1b5cb18732807-1.4-1349388036-0