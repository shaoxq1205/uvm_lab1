/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sce/sce0ae492a37d919f-1.3-1349388176-0