/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s10/s10c0c5fdc6f3976c-1.4-1349388027-0