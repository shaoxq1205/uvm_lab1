/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sb4/sb4d8c24a6a733ad1-1.4-1349388116-0