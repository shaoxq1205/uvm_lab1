/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sd7/sd74024357de6fc9a-1.4-1349388236-0