library verilog;
use verilog.vl_types.all;
entity GlobalPipeInfo is
end GlobalPipeInfo;
