/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s77/s77c62cb6e6ea21b4-1.4-1349388128-0