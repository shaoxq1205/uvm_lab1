/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s99/s998990abd0b1f264-1.4-1349387984-0