/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/se3/se38e9c1a6c2908ba-1.4-1349388132-0