/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s01/s01763ea8ff5f9dfa-1.4-1349388122-0