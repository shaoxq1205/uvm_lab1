/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s44/s44c5e2c33d70bbec-1.4-1349388073-0