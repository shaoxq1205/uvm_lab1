/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s83/s8364f60178641dba-1.4-1349388126-0