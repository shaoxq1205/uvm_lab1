/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s5e/s5e605b480d6848c4-1.4-1349388187-0