library verilog;
use verilog.vl_types.all;
entity XlClockAdvancer is
    port(
        clock           : in     vl_logic
    );
end XlClockAdvancer;
