/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sb1/sb18a6b20d65ff7e0-1.4-1349388135-0