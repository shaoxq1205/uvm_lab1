/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sf9/sf9880945190fa0ab-1.4-1349388195-0