/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sff/sff14a6fc1f5addac-1.4-1349388227-0