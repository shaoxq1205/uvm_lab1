/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s0e/s0e509cefcc13cabf-1.3-1349388099-0