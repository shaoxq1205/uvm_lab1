/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sdf/sdf3ee18971fe3e99-1.4-1349388038-0