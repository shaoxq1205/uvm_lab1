/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/saa/saa9d17984a3aa256-1.4-1349388231-0