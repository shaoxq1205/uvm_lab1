/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s58/s58d164225c59b551-1.4-1349388224-0