library verilog;
use verilog.vl_types.all;
entity XlSvGpioTransactorPkg is
end XlSvGpioTransactorPkg;
