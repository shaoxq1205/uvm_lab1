/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/scb/scbac693c3257bc78-1.4-1349388185-0