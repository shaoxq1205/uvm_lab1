/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s2a/s2a1210663a6f5167-1.3-1349388149-0