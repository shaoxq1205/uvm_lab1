/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s25/s25ff7869aed9b9d3-1.3-1349388173-0