/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s54/s546dd64201d7bcc7-1.4-1349388077-0