/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sf5/sf517d32177a10629-1.4-1349388184-0