/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s9a/s9af5e509d10e7399-1.3-1349388187-0