/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s49/s4945afdfde8858bb-1.4-1349388182-0