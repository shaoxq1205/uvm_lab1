/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sc0/sc0bbdc3e251cc2ba-1.4-1349388187-0