/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s24/s24f9ffb29ff7f563-1.4-1349388117-0