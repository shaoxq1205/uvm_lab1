library verilog;
use verilog.vl_types.all;
entity XlSvTimeAdvancerPkg is
end XlSvTimeAdvancerPkg;
