/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s93/s9374feea65cec491-1.4-1349388194-0