/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sf0/sf0530187ddc57497-1.4-1349387984-0