library verilog;
use verilog.vl_types.all;
entity TbxScManager is
end TbxScManager;
