/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sd6/sd60d8c57549c844d-1.4-1349388092-0