/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s6e/s6eddb443a17860bb-1.4-1349388177-0