/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s6a/s6acc37a6e337c452-1.3-1349388130-0