/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sd0/sd0a8d2216748f7a7-1.4-1349387981-0