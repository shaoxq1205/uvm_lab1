/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s46/s4672ba6c978bb2f6-1.3-1349388186-0