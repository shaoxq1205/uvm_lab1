/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s10/s10ab62d3a62ece07-1.4-1349388235-0