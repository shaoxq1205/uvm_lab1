/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s69/s69025399b6086558-1.4-1349388136-0