library verilog;
use verilog.vl_types.all;
entity XlSvEdgeDetectorPkg is
end XlSvEdgeDetectorPkg;
