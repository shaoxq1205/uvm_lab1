/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sf5/sf53445576fcfeb0b-1.4-1349388134-0