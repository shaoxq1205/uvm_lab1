library verilog;
use verilog.vl_types.all;
entity pcounter_pkg is
end pcounter_pkg;
