/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s33/s331986ce9fb37402-1.3-1349388099-0