/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sc6/sc63fb39e14ff49b3-1.4-1349388219-0