/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sb5/sb50230bb0c265fdb-1.4-1349387983-0