/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s68/s6858693d534846e7-1.4-1349388230-0