/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s27/s2769d5a0e867e233-1.4-1349388179-0