/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s43/s436f19493e14f863-1.4-1349388124-0