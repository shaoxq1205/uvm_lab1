/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s0f/s0fb26dd22326eed5-1.4-1349388196-0