/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s0b/s0b8e727812e6ab30-1.4-1349388020-0