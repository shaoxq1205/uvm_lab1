/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s22/s2269e80f6b8d5fd8-1.4-1349388122-0