/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sa4/sa4f74ce4754758ac-1.4-1349388074-0