package XlSvPkg2;

    `include "XlSvClockAdvancer.svh"
    `include "XlSvResetGenerator.svh"

  
endpackage : XlSvPkg2
