/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sc7/sc783353de28ba871-1.4-1349388195-0