/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s8f/s8f11ea9d4ff276cd-1.4-1349388228-0