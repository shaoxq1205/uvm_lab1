/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sfa/sfaed4bb0f4ba2d3c-1.4-1349388000-0