/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s8d/s8d923ddcea435770-1.4-1349388130-0