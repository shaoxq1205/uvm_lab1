/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s8b/s8b9ac111bf7d401d-1.4-1349388227-0