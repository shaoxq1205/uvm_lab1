/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s72/s72b81d53624a9147-1.4-1349388234-0