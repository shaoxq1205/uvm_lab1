/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sb5/sb51b5392d8132e66-1.4-1349388024-0