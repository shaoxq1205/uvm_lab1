/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s58/s58221358e9ce4468-1.4-1349388001-0