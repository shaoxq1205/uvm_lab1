/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sd6/sd68d56e619ab891a-1.3-1349388148-0