/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s64/s64e0fa75fb5e0266-1.4-1349387983-0