/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s9b/s9b56e638fa9f0df9-1.4-1349388003-0