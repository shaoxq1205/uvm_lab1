/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/se0/se022c5b6d314098d-1.4-1349388017-0