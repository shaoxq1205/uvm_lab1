/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sbf/sbfc69f084435c190-1.4-1349388141-0