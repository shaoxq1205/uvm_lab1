/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sfe/sfee075cabf12c56b-1.4-1349387969-0