/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s8c/s8c363b8224713186-1.4-1349388224-0