/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s7a/s7af209868ae018cd-1.4-1349388231-0