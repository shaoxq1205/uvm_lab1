/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s0f/s0f3250b12fb0a1b6-1.4-1349388234-0