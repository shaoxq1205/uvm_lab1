/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s68/s6887af2421dc0015-1.3-1349388099-0