/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s29/s2938ca916f8e0ac3-1.4-1349388176-0