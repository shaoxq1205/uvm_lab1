/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s2a/s2aaf6ae62fca3f41-1.4-1349388012-0