/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s7c/s7c27c2fda3b3c454-1.4-1349388121-0