/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s07/s07c877c2f26d1e0b-1.4-1349388127-0