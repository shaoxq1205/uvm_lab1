/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/se2/se29ca44e5829578c-1.4-1349388119-0