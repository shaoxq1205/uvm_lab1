/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sff/sff7c6d43b25e0a2b-1.4-1349388186-0