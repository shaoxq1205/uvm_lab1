/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/saa/saab966b7c633ba9f-1.4-1349388137-0