/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/scb/scb46084392dad9ce-1.4-1349388017-0