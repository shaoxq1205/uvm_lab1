/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s7b/s7bccfc4d301944b5-1.4-1349388027-0