/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/se3/se366bbf04851e677-1.4-1349388008-0