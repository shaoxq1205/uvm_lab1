/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s29/s29db6a108f33ba98-1.4-1349388119-0