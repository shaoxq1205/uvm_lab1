/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s9c/s9c784bc86001f51d-1.4-1349388141-0