/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s17/s1791894cd4439e33-1.4-1349388003-0