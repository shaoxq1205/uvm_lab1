/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sdd/sddaecdee98a5b45c-1.3-1349388016-0