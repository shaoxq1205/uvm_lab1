/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sfd/sfd9d9f15bcc63089-1.4-1349388016-0