/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s75/s7579401cb29889e9-1.4-1349388123-0