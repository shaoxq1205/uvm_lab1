/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s02/s023e0c3b832190e6-1.4-1349388021-0