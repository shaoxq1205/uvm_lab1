/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s86/s86a036a5a68cd5d1-1.4-1349388181-0