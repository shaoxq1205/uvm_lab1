/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sbe/sbe43a517d0b430c9-1.4-1349388019-0