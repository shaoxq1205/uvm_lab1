/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s54/s54f0d10e18160827-1.4-1349388133-0