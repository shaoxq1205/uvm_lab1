/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s03/s038e661271a477d5-1.4-1349388155-0