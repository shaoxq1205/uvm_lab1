/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sf9/sf93334db1e1fb26c-1.4-1349388192-0