/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/seb/seb22d581fd5bb467-1.4-1349388028-0