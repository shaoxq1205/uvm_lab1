/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s8a/s8a373f3f2799da03-1.4-1349387982-0