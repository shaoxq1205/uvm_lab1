library verilog;
use verilog.vl_types.all;
entity XlVeraSystemClock is
    port(
        clock           : in     vl_logic
    );
end XlVeraSystemClock;
