/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s26/s26f6a71b43d60048-1.4-1349388125-0