/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sed/sedca52bd36fb0b12-1.4-1349388226-0