/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sa9/sa969dfef08901373-1.3-1349388149-0