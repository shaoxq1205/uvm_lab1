/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sd4/sd4c33674f472dd9f-1.4-1349388189-0