/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s4b/s4b7254035fba6d71-1.4-1349388039-0