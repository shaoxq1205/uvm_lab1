/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sd8/sd82c1ab36faac0b0-1.4-1349388177-0