/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s2d/s2d15a555043f8d99-1.4-1349388191-0