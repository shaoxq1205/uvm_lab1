//-----------------------------------------------------------------------------
// Qualcomm Proprietary
// Copyright (c) Qualcomm Inc.
// All rights reserved.
//
//
// All data and information contained in or disclosed by this document
// are confidential and proprietary information of QUALCOMM Incorporated,
// and all rights therein are expressly reserved. By accepting this
// material, the recipient agrees that this material and the information
// contained therein are held in confidence and in trust and will not be
// used, copied, reproduced in whole or in part, nor its contents
// revealed in any manner to others without the express written
// permission of QUALCOMM Incorporated.
//
// This technology was exported from the United States in accordance with
// the Export Administration Regulations. Diversion contrary to U.S. law
// prohibited.
//-----------------------------------------------------------------------------
/**
 * @brief Pcounter Sequence List
 *
 * The Pcounter DUT Sequence List File (pcounter_seq_list.sv) contains all 
 * of the available sequences for the Pcounter DUT.
 *
 * @file pcounter_seq_list.sv
 *
 * @author Loganath Ramachandran
 * @par Contact:
 * c_lramc@qualcomm.com
 * @par Location:
 * QC-SD
 *
 * $Revision: 1.3 $
 * $Date: Mon Nov 15 12:05:24 2010 $
 * $Author: mironm $
 */

`ifndef PCOUNTER_SEQ_LIST__SV
`define PCOUNTER_SEQ_LIST__SV

`include "uvm_macros.svh"
import uvm_pkg::*;


`include "pcounter_test_qclk_change_clock_period_vseq.sv"


`endif
