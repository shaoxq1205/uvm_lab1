/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s62/s626073cf5d9385e2-1.4-1349388195-0