/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s9d/s9de84dbd51e0d10a-1.4-1349388026-0