/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s46/s467f60f5123ad444-1.4-1349388093-0