/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s69/s69437773ac3d7cfe-1.4-1349388139-0