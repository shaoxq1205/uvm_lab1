/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s1b/s1b69542ed439cd87-1.4-1349388151-0