/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sd3/sd3683146a9f1594b-1.4-1349387995-0