/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sce/sce0e7fe426283823-1.4-1349388157-0