/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sa9/sa973812d4f13efe4-1.3-1349388124-0