/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s00/s00324155e7fae9c9-1.4-1349388121-0