/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/scb/scb1b25fb93368dfa-1.4-1349387997-0