/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sb4/sb41964e947ee9ffd-1.4-1349388189-0