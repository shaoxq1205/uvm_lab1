/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s3b/s3b66c93432f341c3-1.4-1349388076-0