/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s98/s98d71905b1f2319f-1.4-1349388199-0