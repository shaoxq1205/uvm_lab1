/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s7d/s7d51c53963bf729d-1.4-1349387967-0