/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/se1/se110714cd18fd39f-1.4-1349388140-0