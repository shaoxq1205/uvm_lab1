library verilog;
use verilog.vl_types.all;
entity XlSvMemoryTransactorPkg is
end XlSvMemoryTransactorPkg;
