/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s1d/s1dfed7f6edf33d02-1.4-1349388152-0