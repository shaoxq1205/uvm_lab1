/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s61/s61bdf1757cf3a810-1.4-1349388172-0