/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sb8/sb8327661b8d31350-1.4-1349388077-0