/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sa4/sa49d67f4ad3caaa1-1.4-1349388224-0