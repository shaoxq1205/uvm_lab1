/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sd5/sd5a6794782dde409-1.4-1349388019-0