/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s37/s377dcab2557d0cbd-1.4-1349388155-0