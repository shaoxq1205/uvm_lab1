/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s6a/s6af08ad02c9cdcef-1.4-1349387995-0