/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s4e/s4e7c5dd11f6c3ca9-1.4-1349387967-0