/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s35/s35d4c14c85e402c0-1.4-1349388180-0