/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s1f/s1fab7720ca0288aa-1.4-1349388128-0