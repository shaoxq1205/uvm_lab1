/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s74/s7446b56b64d226cf-1.4-1349388135-0