library verilog;
use verilog.vl_types.all;
entity xtlm_pkg is
end xtlm_pkg;
