/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sfe/sfea84aeba91fe39b-1.4-1349387988-0