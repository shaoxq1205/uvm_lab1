/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sa8/sa81b125a6e513725-1.4-1349388180-0