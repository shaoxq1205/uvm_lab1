/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sca/sca9f67517f90dcf7-1.4-1349388137-0