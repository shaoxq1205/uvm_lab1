/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s7d/s7dc60d214c8e16d5-1.3-1349388131-0