/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s42/s428bbe846fd65507-1.1-1300484079-0