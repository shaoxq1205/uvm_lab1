/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s64/s64a318ad66ece6a7-1.4-1349388117-0