/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s4b/s4bdff059f97f8580-1.4-1349388010-0