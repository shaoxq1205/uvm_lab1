/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s62/s62901d1fe2c7d6f0-1.4-1349388141-0