/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s19/s19d50a921ea045ad-1.4-1349388222-0