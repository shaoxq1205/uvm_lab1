/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s1a/s1a18ab0c2ae5e02e-1.4-1349388175-0