/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sab/sabd14dee25a09674-1.4-1349388137-0