/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sd6/sd682896f991ffd56-1.4-1349388037-0