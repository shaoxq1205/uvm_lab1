/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s5a/s5a760103b4e37875-1.4-1349388027-0