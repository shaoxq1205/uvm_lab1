/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sa0/sa08992a155be7497-1.4-1349388091-0