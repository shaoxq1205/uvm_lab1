/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sa9/sa9c810a6b7e63eba-1.4-1349388130-0