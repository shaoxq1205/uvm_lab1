/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sa5/sa582c398c1dc825b-1.4-1349388008-0