library verilog;
use verilog.vl_types.all;
entity vsms5505 is
    generic(
        DATA_WIDTH      : integer := 64;
        ID_WIDTH        : integer := 4;
        FIFO_DEPTH      : integer := 8;
        p_resp          : integer := 0;
        p_ch1_id        : integer := 33;
        p_ch2_id        : integer := 34;
        p_ch3_id        : integer := 65;
        p_ch4_id        : integer := 66;
        p_ch1_mask      : integer := 31;
        p_ch2_mask      : integer := 31;
        p_ch3_mask      : integer := 31;
        p_ch4_mask      : integer := 31
    );
    port(
        aclk            : in     vl_logic;
        aresetn         : in     vl_logic;
        arreadyNumWaits_fire: in     vl_logic;
        awreadyNumWaits_fire: in     vl_logic;
        wreadyNumWaits_fire: in     vl_logic;
        awid_p1         : in     vl_logic_vector;
        awaddr_p1       : in     vl_logic_vector(31 downto 0);
        awlen_p1        : in     vl_logic_vector(3 downto 0);
        awsize_p1       : in     vl_logic_vector(2 downto 0);
        awburst_p1      : in     vl_logic_vector(1 downto 0);
        awlock_p1       : in     vl_logic_vector(1 downto 0);
        awcache_p1      : in     vl_logic_vector(3 downto 0);
        awprot_p1       : in     vl_logic_vector(2 downto 0);
        awvalid_p1      : in     vl_logic;
        awready_p1      : out    vl_logic;
        wid_p1          : in     vl_logic_vector;
        wdata_p1        : in     vl_logic_vector;
        wstrb_p1        : in     vl_logic_vector;
        wlast_p1        : in     vl_logic;
        wvalid_p1       : in     vl_logic;
        wready_p1       : out    vl_logic;
        bid_p1          : out    vl_logic_vector;
        bresp_p1        : out    vl_logic_vector(1 downto 0);
        bvalid_p1       : out    vl_logic;
        bready_p1       : in     vl_logic;
        arid_p1         : in     vl_logic_vector;
        araddr_p1       : in     vl_logic_vector(31 downto 0);
        arlen_p1        : in     vl_logic_vector(3 downto 0);
        arsize_p1       : in     vl_logic_vector(2 downto 0);
        arburst_p1      : in     vl_logic_vector(1 downto 0);
        arlock_p1       : in     vl_logic_vector(1 downto 0);
        arcache_p1      : in     vl_logic_vector(3 downto 0);
        arprot_p1       : in     vl_logic_vector(2 downto 0);
        arvalid_p1      : in     vl_logic;
        arready_p1      : out    vl_logic;
        rid_p1          : out    vl_logic_vector;
        rdata_p1        : out    vl_logic_vector;
        rresp_p1        : out    vl_logic_vector(1 downto 0);
        rlast_p1        : out    vl_logic;
        rvalid_p1       : out    vl_logic;
        rready_p1       : in     vl_logic;
        awid_p2         : in     vl_logic_vector;
        awaddr_p2       : in     vl_logic_vector(31 downto 0);
        awlen_p2        : in     vl_logic_vector(3 downto 0);
        awsize_p2       : in     vl_logic_vector(2 downto 0);
        awburst_p2      : in     vl_logic_vector(1 downto 0);
        awlock_p2       : in     vl_logic_vector(1 downto 0);
        awcache_p2      : in     vl_logic_vector(3 downto 0);
        awprot_p2       : in     vl_logic_vector(2 downto 0);
        awvalid_p2      : in     vl_logic;
        awready_p2      : out    vl_logic;
        wid_p2          : in     vl_logic_vector;
        wdata_p2        : in     vl_logic_vector;
        wstrb_p2        : in     vl_logic_vector;
        wlast_p2        : in     vl_logic;
        wvalid_p2       : in     vl_logic;
        wready_p2       : out    vl_logic;
        bid_p2          : out    vl_logic_vector;
        bresp_p2        : out    vl_logic_vector(1 downto 0);
        bvalid_p2       : out    vl_logic;
        bready_p2       : in     vl_logic;
        arid_p2         : in     vl_logic_vector;
        araddr_p2       : in     vl_logic_vector(31 downto 0);
        arlen_p2        : in     vl_logic_vector(3 downto 0);
        arsize_p2       : in     vl_logic_vector(2 downto 0);
        arburst_p2      : in     vl_logic_vector(1 downto 0);
        arlock_p2       : in     vl_logic_vector(1 downto 0);
        arcache_p2      : in     vl_logic_vector(3 downto 0);
        arprot_p2       : in     vl_logic_vector(2 downto 0);
        arvalid_p2      : in     vl_logic;
        arready_p2      : out    vl_logic;
        rid_p2          : out    vl_logic_vector;
        rdata_p2        : out    vl_logic_vector;
        rresp_p2        : out    vl_logic_vector(1 downto 0);
        rlast_p2        : out    vl_logic;
        rvalid_p2       : out    vl_logic;
        rready_p2       : in     vl_logic;
        csysreq         : in     vl_logic;
        csysack         : in     vl_logic;
        cactive         : in     vl_logic;
        i_sram_d        : in     vl_logic_vector;
        o_sram_q        : out    vl_logic_vector;
        o_sram_waddr    : out    vl_logic_vector(31 downto 0);
        o_sram_raddr    : out    vl_logic_vector(31 downto 0);
        o_sram_be       : out    vl_logic_vector(15 downto 0);
        o_sram_we       : out    vl_logic;
        o_sram_cs       : out    vl_logic;
        o_sram_clk      : out    vl_logic
    );
end vsms5505;
