/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/scc/sccd9949656f37932-1.4-1349387982-0