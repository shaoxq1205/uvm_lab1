/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s53/s5323da6cb5108090-1.4-1349388199-0