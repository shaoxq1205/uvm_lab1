/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/scd/scdca312b47f56bea-1.4-1349387988-0