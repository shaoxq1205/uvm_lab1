/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s96/s965276e73ae8adf2-1.4-1349388006-0