/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s1b/s1bd5880465a40740-1.4-1349387989-0