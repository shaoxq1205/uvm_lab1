/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s29/s298436054c972642-1.4-1349388192-0