/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s0a/s0aabe087a6435675-1.4-1349388038-0