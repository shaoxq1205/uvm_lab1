/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s91/s91f4f941ad854e4b-1.4-1349388183-0