/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s74/s745c7cc22ad744cb-1.4-1349388091-0