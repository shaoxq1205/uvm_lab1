/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s33/s33b76f5c82b597ed-1.4-1349388151-0