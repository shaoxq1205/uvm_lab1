/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sb4/sb403c99941b887b3-1.4-1349388190-0