/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sc5/sc55f369339c93a32-1.4-1349388190-0