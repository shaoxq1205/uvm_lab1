/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s39/s39843374a759358c-1.4-1349388191-0