/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s9b/s9bf16d5bba367158-1.4-1349388156-0