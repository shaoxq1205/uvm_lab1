/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s9b/s9b28f3d189001ceb-1.4-1349388005-0