/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s9c/s9c2c0caf5f9dffce-1.4-1349388229-0