library verilog;
use verilog.vl_types.all;
entity XlSvPkg is
end XlSvPkg;
