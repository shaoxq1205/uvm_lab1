/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sfc/sfcfa9ad32860d71a-1.4-1349388129-0