/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sc3/sc3fca4968ddb6b91-1.4-1349388129-0