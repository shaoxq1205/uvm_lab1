/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sf5/sf5863539e864c708-1.3-1349388147-0