/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sbd/sbdadfde1426ec09d-1.4-1349388025-0