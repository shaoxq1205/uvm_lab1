/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s2b/s2beca7de119dbf71-1.4-1349388198-0