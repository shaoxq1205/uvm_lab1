/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sb9/sb9a89310f16a227c-1.4-1349388182-0