/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sa4/sa40caf9a63d2d4a7-1.4-1349388017-0