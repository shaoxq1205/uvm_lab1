/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s1a/s1a413d5f68278130-1.4-1349388004-0