/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sdc/sdc7152176af18ec8-1.4-1349388156-0