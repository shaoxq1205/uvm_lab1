/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sca/scac4b327cc490665-1.3-1349388071-0