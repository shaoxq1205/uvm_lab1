/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sb0/sb02ec30ad562904e-1.4-1349388008-0