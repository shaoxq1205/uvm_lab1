/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sba/sbada614491cf0e81-1.4-1349387970-0