/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s23/s23a280a9542df604-1.4-1349388196-0