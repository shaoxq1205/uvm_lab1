/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sa6/sa6f85fb0be24c982-1.4-1349388018-0