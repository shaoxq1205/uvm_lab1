/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s06/s0619cff2b8d21d36-1.4-1349388179-0