/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sb7/sb7af08b8eba4b2db-1.3-1349388002-0