/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sa5/sa5103391f2be5cd4-1.4-1349388132-0