/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/se9/se915ad57db88bf9a-1.4-1349388174-0