/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s70/s70f3a5dbb1c9d1cb-1.4-1349388235-0