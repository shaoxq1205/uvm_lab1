/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s22/s22cfad52c7342a5e-1.4-1349388159-0