/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s1d/s1daa404c8e6c1dfa-1.4-1349387997-0