/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/se4/se478714bdad91ab4-1.4-1349388179-0