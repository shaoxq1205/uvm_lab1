/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sc0/sc03987a764e0f62e-1.3-1349388098-0