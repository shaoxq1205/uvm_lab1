/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sed/sedcc189ade31dafd-1.4-1349388142-0