library verilog;
use verilog.vl_types.all;
entity tbx_event_pkg is
end tbx_event_pkg;
