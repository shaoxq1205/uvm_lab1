/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sd5/sd564c1e79a946368-1.4-1349388123-0