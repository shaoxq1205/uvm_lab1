/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s67/s67fb22e291f6f92b-1.4-1349388131-0