/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sd7/sd77103b65bbd5fd4-1.4-1349387985-0