/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/scf/scf858dc30e90f160-1.3-1349388071-0