/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s2b/s2b940b733e78d3b4-1.4-1349388181-0