/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s16/s167537dbd5ae0640-1.4-1349388220-0