/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s3d/s3d8dc862d5c76ffe-1.4-1349388193-0