/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sa1/sa136f14210b42362-1.3-1349388174-0