/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sb7/sb785e755f9c06a6e-1.4-1349388124-0