/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sf3/sf3e6097db0f84450-1.4-1349388183-0