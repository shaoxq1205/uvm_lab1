/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sbf/sbfb08b76ed4deb87-1.3-1349388147-0