/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s1e/s1eb0a352f431ed66-1.4-1349388175-0