/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/se2/se2209505fa038a91-1.4-1349388120-0