/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s6b/s6b4bb6622d2ec735-1.4-1349388039-0