/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s18/s188845a3e717383c-1.4-1349388173-0