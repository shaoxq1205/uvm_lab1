/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sa1/sa168ec23350a7418-1.4-1349388022-0