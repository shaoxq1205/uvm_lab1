/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s7c/s7c12e00e986ef996-1.4-1349388010-0