/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/scd/scd26774c928e5bf9-1.4-1349388093-0