/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s94/s94a61284d6f9c0cf-1.4-1349388125-0