/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s3b/s3bac0b5b41edd13f-1.4-1349388194-0