/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/se1/se162b49cc441531a-1.4-1349388194-0