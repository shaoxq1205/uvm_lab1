/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sad/sad533eed21263072-1.4-1349388089-0