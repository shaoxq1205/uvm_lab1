/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s28/s288ee18580ee9d59-1.4-1349388236-0