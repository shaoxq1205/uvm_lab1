/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s44/s4454c6a9e7dbeeee-1.4-1349388091-0