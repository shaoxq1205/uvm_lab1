/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sf8/sf8bbd14007a2dfd5-1.4-1349388136-0