/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s5a/s5ada4e76b52e14bb-1.4-1349388158-0