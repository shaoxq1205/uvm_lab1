/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s72/s7224a8a03e1ab67a-1.4-1349388117-0