/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s11/s114bdd5b7e18e27a-1.4-1349388197-0