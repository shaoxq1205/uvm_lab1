/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s30/s3037c2f85647f28a-1.4-1349388073-0