/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sdf/sdf025b1237d33cec-1.4-1349388018-0