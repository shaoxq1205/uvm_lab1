/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sb4/sb4edd06b3cba6dd4-1.4-1349388010-0