/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s00/s007ecb565f369a40-1.4-1349388191-0