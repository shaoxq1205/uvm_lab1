/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s56/s5633b0917ac58d01-1.4-1349388001-0