/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s2b/s2b7105c94744960e-1.4-1349388004-0