/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s05/s053dc16d74c25c65-1.4-1349388221-0