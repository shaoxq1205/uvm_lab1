library verilog;
use verilog.vl_types.all;
entity qclk_pkg is
end qclk_pkg;
