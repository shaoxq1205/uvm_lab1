/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s02/s025a53dbd096b0df-1.4-1349388074-0