/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sec/sec59efcffbb483df-1.4-1349388153-0