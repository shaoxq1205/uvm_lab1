/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s63/s636644472d56f8d9-1.4-1349388076-0