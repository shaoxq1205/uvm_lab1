/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s49/s4993f0526c03a214-1.4-1349387983-0