/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sf5/sf59a4dd3749dfb6c-1.4-1349387987-0