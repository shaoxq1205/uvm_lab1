/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s0a/s0aaa74407e4eb5df-1.4-1349388189-0