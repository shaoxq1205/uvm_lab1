/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s72/s728e5f357f4913c6-1.4-1349388134-0