/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s9a/s9abcd7be9f7ab06c-1.4-1349388024-0