/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s8f/s8f771d52aebddcbb-1.4-1349388235-0