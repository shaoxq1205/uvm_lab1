/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sc2/sc2f80d9981a62b56-1.4-1349387996-0