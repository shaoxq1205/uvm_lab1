/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s23/s23e30167931c29cd-1.4-1349388178-0