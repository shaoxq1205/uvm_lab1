/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s36/s36359ad94c23ac88-1.4-1349388156-0