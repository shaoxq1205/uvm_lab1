/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sde/sde6ae3437b7f306d-1.2-1350508795-0