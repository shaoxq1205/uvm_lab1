/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s70/s70ac98c7056c05c7-1.4-1349388073-0