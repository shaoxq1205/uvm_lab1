/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s67/s67d6d266cc02bd9e-1.4-1349388089-0