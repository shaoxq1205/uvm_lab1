/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sc8/sc83bb1039edf355c-1.4-1349388005-0