/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s63/s632cd315b42f3a48-1.4-1349388128-0