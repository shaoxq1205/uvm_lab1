/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s19/s198642309607c6a7-1.3-1349388173-0