/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s81/s81a48d6bfdfbf051-1.4-1349387985-0