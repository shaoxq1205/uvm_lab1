/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s4a/s4a6b8bd3aa631148-1.4-1349388185-0