/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sca/scad00caec55218ab-1.4-1349387984-0