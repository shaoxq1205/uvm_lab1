/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/se1/se137cbaf1dff1f80-1.4-1349388000-0