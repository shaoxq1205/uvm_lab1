/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s8d/s8d9551a19da8153b-1.4-1349388011-0