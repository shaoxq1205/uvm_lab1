/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s5d/s5dbbde7d56c09e64-1.4-1349388196-0