/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sf2/sf2cc1fed12a7c913-1.4-1349387996-0