library verilog;
use verilog.vl_types.all;
entity xtlm_base_pkg is
end xtlm_base_pkg;
