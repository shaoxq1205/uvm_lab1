/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s13/s1359f1b5d24b1874-1.4-1349388159-0