/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s6c/s6c2e27638a546236-1.4-1349388000-0