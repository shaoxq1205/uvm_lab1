/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/se9/se931d628020474a2-1.4-1349388003-0