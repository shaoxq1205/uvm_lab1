/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s1a/s1a57ca5852a3aea1-1.4-1349387997-0