/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s92/s922ee5518e7217f2-1.4-1349388002-0