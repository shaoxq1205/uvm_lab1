/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s62/s6253f8c9b599398b-1.4-1349388011-0