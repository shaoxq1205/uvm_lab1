library verilog;
use verilog.vl_types.all;
entity tbx_internal_DumpExport_Defns_SIM is
end tbx_internal_DumpExport_Defns_SIM;
