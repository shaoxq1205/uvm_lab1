/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s9b/s9b8b00d098e1259c-1.4-1349388226-0