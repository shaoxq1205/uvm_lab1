library verilog;
use verilog.vl_types.all;
entity TbxSvManager is
end TbxSvManager;
