/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s56/s56ad9e6d7eae67a2-1.4-1349388130-0