/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s31/s3112472c198f85b1-1.4-1349388151-0