/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s43/s43a7a21c33dc530b-1.4-1349388185-0