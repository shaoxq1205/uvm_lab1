/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s4f/s4f808e05d522cebd-1.4-1349388183-0