/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/see/see69dc4e927d0cf8-1.4-1349388134-0