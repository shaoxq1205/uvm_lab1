/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s5b/s5bf3d03fa50c9a9f-1.4-1349388220-0