/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s40/s4031624619e38abb-1.3-1349388186-0