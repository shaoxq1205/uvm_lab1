/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sb7/sb7abe0975698a0eb-1.4-1349388158-0