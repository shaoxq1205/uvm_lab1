/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s25/s25d64487b960f3ee-1.4-1349388178-0