/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sef/sef0a5d158e95ddf0-1.4-1349388013-0