/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s6c/s6cab44d1702bf948-1.4-1349388232-0