/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sd7/sd74b1a7a598d47bb-1.4-1349388158-0