/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s34/s34e40673560fc117-1.4-1349387967-0