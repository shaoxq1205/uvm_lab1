/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s38/s38e8fffa60e99c4b-1.4-1349388160-0