/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/s1c/s1ce45bb3eae163c2-1.4-1349388197-0