/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sa9/sa97b80c1bc20a1bc-1.4-1349388074-0