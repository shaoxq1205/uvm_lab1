/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/se9/se94db7e405915194-1.4-1349388155-0