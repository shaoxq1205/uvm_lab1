/prj/qct/verif/svtb/sandiego/.synchronicity/sync_cache/sfd/sfdc61ed2d37cabeb-1.4-1349388037-0